module riscv_imm_gen(

) (

)

endmodule
